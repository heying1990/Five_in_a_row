library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity table_fifteen is
    Port (Reset : in std_logic;
          frame_clk : in std_logic;
          state_out : in std_logic_vector(3 downto 0);
          Button : in std_logic_vector(7 downto 0);
          block00X : out std_logic_vector(9 downto 0);
          block00Y : out std_logic_vector(9 downto 0);
          block01X : out std_logic_vector(9 downto 0);
          block01Y : out std_logic_vector(9 downto 0);
          block02X : out std_logic_vector(9 downto 0);
          block02Y : out std_logic_vector(9 downto 0);
          block03X : out std_logic_vector(9 downto 0);
          block03Y : out std_logic_vector(9 downto 0);
          block04X : out std_logic_vector(9 downto 0);
          block04Y : out std_logic_vector(9 downto 0);
          block05X : out std_logic_vector(9 downto 0);
          block05Y : out std_logic_vector(9 downto 0);
          
          
          chess_positionX : out std_logic_vector(9 downto 0);
          chess_positionY : out std_logic_vector(9 downto 0);
          chess_size : out std_logic_vector(9 downto 0);
          stopsig : out std_logic);

end table_fifteen;

architecture Behavioral of table_fifteen is
signal movingX : std_logic_vector(9 downto 0);
signal movingY : std_logic_vector(9 downto 0);
signal chess_motionX : std_logic_vector(9 downto 0);
signal chess_motionY : std_logic_vector(9 downto 0);
signal counter : std_logic_vector(9 downto 0);
signal stop : std_logic;
signal size : std_logic_vector(9 downto 0);

constant chess_centerX : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 335,10);
constant chess_centerY : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 255,10);
constant chess_stepX : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(2 ,10);
constant chess_stepY : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(2 ,10);

constant chess_maxX :  std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 555,10);
constant chess_maxY :  std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 475,10);
constant chess_minX :  std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 115,10);
constant chess_minY :  std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 35,10);

constant chess_centerX : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 335,10);
constant chess_centerY : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 255,10);
constant chess_stepX : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(2 ,10);
constant chess_stepY : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(2 ,10);

constant block00X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(125,10);
constant block00Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 45,10);
constant block01X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 155,10);
constant block01Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 45,10);
constant block02X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 185,10);
constant block02Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 45,10);
constant block03X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 215,10);
constant block03Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 45,10);
constant block04X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 245,10);
constant block04Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 45,10);
constant block05X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 275,10);
constant block05Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 45,10);
constant block06X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 305,10);
constant block06Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 45,10);
constant block07X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 335,10);
constant block07Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 45,10);
constant block08X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 365,10);
constant block08Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 45,10);
constant block09X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 395,10);
constant block09Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 45,10);
constant block10X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 425,10);
constant block10Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 45,10);
constant block11X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 455,10);
constant block11Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 45,10);
constant block12X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 485,10);
constant block12Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 45,10);
constant block13X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 515,10);
constant block13Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 45,10);
constant block14X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 545,10);
constant block14Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 45,10);
constant block15X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(125,10);
constant block15Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 75,10);
constant block16X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 155,10);
constant block16Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 75,10);
constant block17X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 185,10);
constant block17Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 75,10);
constant block18X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 215,10);
constant block18Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 75,10);
constant block19X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 245,10);
constant block19Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 75,10);
constant block20X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 275,10);
constant block20Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 75,10);
constant block21X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 305,10);
constant block21Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 75,10);
constant block22X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 335,10);
constant block22Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 75,10);
constant block23X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 365,10);
constant block23Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 75,10);
constant block24X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 395,10);
constant block24Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 75,10);
constant block25X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 425,10);
constant block25Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 75,10);
constant block26X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 455,10);
constant block26Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 75,10);
constant block27X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 485,10);
constant block27Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 75,10);
constant block28X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 515,10);
constant block28Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 75,10);
constant block29X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 545,10);
constant block29Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 75,10);
constant block30X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR(125,10);
constant block30Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 105,10);
constant block31X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 155,10);
constant block31Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 105,10);
constant block32X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 185,10);
constant block32Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 105,10);
constant block33X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 215,10);
constant block33Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 105,10);
constant block34X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 245,10);
constant block34Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 105,10);
constant block35X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 275,10);
constant block35Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 105,10);
constant block36X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 305,10);
constant block36Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 105,10);
constant block37X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 335,10);
constant block37Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 105,10);
constant block38X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 365,10);
constant block38Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 105,10);
constant block39X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 395,10);
constant block39Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 105,10);
constant block40X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 425,10);
constant block40Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 105,10);
constant block41X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 455,10);
constant block41Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 105,10);
constant block42X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 485,10);
constant block42Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 105,10);
constant block43X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 515,10);
constant block43Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 105,10);
constant block44X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 545,10);
constant block44Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 105,10);
constant block45X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 125,10);
constant block45Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 135,10);
constant block46X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 155,10);
constant block46Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 135,10);
constant block47X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 185,10);
constant block47Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 135,10);
constant block48X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 215,10);
constant block48Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 135,10);
constant block49X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 245,10);
constant block49Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 135,10);
constant block50X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 275,10);
constant block50Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 135,10);
constant block51X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 305,10);
constant block51Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 135,10);
constant block52X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 335,10);
constant block52Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 135,10);
constant block53X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 365,10);
constant block53Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 135,10);
constant block54X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 395,10);
constant block54Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 135,10);
constant block55X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 425,10);
constant block55Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 135,10);
constant block56X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 455,10);
constant block56Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 135,10);
constant block57X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 485,10);
constant block57Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 135,10);
constant block58X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 515,10);
constant block58Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 135,10);
constant block59X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 545,10);
constant block59Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 135,10);
constant block60X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 125,10);
constant block60Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 165,10);
constant block61X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 155,10);
constant block61Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 165,10);
constant block62X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 185,10);
constant block62Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 165,10);
constant block63X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 215,10);
constant block63Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 165,10);
constant block64X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 245,10);
constant block64Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 165,10);
constant block65X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 275,10);
constant block65Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 165,10);
constant block66X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 305,10);
constant block66Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 165,10);
constant block67X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 335,10);
constant block67Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 165,10);
constant block68X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 365,10);
constant block68Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 165,10);
constant block69X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 395,10);
constant block69Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 165,10);
constant block70X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 425,10);
constant block70Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 165,10);
constant block71X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 455,10);
constant block71Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 165,10);
constant block72X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 485,10);
constant block72Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 165,10);
constant block73X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 515,10);
constant block73Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 165,10);
constant block74X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 545,10);
constant block74Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 165,10);
constant block75X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 125,10);
constant block75Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 195,10);
constant block76X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 155,10);
constant block76Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 195,10);
constant block77X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 185,10);
constant block77Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 195,10);
constant block78X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 215,10);
constant block78Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 195,10);
constant block79X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 245,10);
constant block79Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 195,10);
constant block80X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 275,10);
constant block80Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 195,10);
constant block81X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 305,10);
constant block81Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 195,10);
constant block82X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 335,10);
constant block82Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 195,10);
constant block83X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 365,10);
constant block83Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 195,10);
constant block84X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 395,10);
constant block84Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 195,10);
constant block85X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 425,10);
constant block85Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 195,10);
constant block86X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 455,10);
constant block86Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 195,10);
constant block87X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 485,10);
constant block87Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 195,10);
constant block88X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 515,10);
constant block88Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 195,10);
constant block89X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 545,10);
constant block89Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 195,10);
constant block90X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 125,10);
constant block90Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 225,10);
constant block91X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 155,10);
constant block91Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 225,10);
constant block92X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 185,10);
constant block92Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 225,10);
constant block93X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 215,10);
constant block93Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 225,10);
constant block94X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 245,10);
constant block94Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 225,10);
constant block95X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 275,10);
constant block95Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 225,10);
constant block96X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 305,10);
constant block96Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 225,10);
constant block97X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 335,10);
constant block97Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 225,10);
constant block98X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 365,10);
constant block98Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 225,10);
constant block99X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 395,10);
constant block99Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 225,10);
constant block100X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 425,10);
constant block100Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 225,10);
constant block101X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 455,10);
constant block101Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 225,10);
constant block102X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 485,10);
constant block102Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 225,10);
constant block103X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 515,10);
constant block103Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 225,10);
constant block104X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 545,10);
constant block104Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 225,10);
constant block105X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 125,10);
constant block105Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 255,10);
constant block106X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 155,10);
constant block106Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 255,10);
constant block107X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 185,10);
constant block107Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 255,10);
constant block108X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 215,10);
constant block108Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 255,10);
constant block109X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 245,10);
constant block109Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 255,10);
constant block110X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 275,10);
constant block110Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 255,10);
constant block111X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 305,10);
constant block111Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 255,10);
constant block112X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 335,10);
constant block112Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 255,10);
constant block113X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 365,10);
constant block113Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 255,10);
constant block114X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 395,10);
constant block114Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 255,10);
constant block115X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 425,10);
constant block115Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 255,10);
constant block116X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 455,10);
constant block116Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 255,10);
constant block117X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 485,10);
constant block117Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 255,10);
constant block118X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 515,10);
constant block118Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 255,10);
constant block119X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 545,10);
constant block119Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 255,10);
constant block120X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 125,10);
constant block120Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 285,10);
constant block121X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 155,10);
constant block121Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 285,10);
constant block122X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 185,10);
constant block122Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 285,10);
constant block123X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 215,10);
constant block123Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 285,10);
constant block124X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 245,10);
constant block124Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 285,10);
constant block125X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 275,10);
constant block125Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 285,10);
constant block126X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 305,10);
constant block126Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 285,10);
constant block127X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 335,10);
constant block127Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 285,10);
constant block128X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 365,10);
constant block128Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 285,10);
constant block129X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 395,10);
constant block129Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 285,10);
constant block130X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 425,10);
constant block130Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 285,10);
constant block131X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 455,10);
constant block131Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 285,10);
constant block132X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 485,10);
constant block132Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 285,10);
constant block133X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 515,10);
constant block133Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 285,10);
constant block134X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 545,10);
constant block134Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 285,10);
constant block135X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 125,10);
constant block135Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 315,10);
constant block136X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 155,10);
constant block136Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 315,10);
constant block137X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 185,10);
constant block137Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 315,10);
constant block138X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 215,10);
constant block138Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 315,10);
constant block139X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 245,10);
constant block139Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 315,10);
constant block140X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 275,10);
constant block140Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 315,10);
constant block141X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 305,10);
constant block141Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 315,10);
constant block142X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 335,10);
constant block142Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 315,10);
constant block143X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 365,10);
constant block143Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 315,10);
constant block144X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 395,10);
constant block144Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 315,10);
constant block145X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 425,10);
constant block145Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 315,10);
constant block146X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 455,10);
constant block146Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 315,10);
constant block147X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 485,10);
constant block147Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 315,10);
constant block148X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 515,10);
constant block148Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 315,10);
constant block149X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 545,10);
constant block149Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 315,10);
constant block150X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 125,10);
constant block150Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 345,10);
constant block151X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 155,10);
constant block151Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 345,10);
constant block152X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 185,10);
constant block152Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 345,10);
constant block153X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 215,10);
constant block153Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 345,10);
constant block154X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 245,10);
constant block154Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 345,10);
constant block155X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 275,10);
constant block155Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 345,10);
constant block156X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 305,10);
constant block156Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 345,10);
constant block157X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 335,10);
constant block157Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 345,10);
constant block158X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 365,10);
constant block158Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 345,10);
constant block159X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 395,10);
constant block159Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 345,10);
constant block160X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 425,10);
constant block160Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 345,10);
constant block161X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 455,10);
constant block161Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 345,10);
constant block162X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 485,10);
constant block162Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 345,10);
constant block163X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 515,10);
constant block163Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 345,10);
constant block164X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 545,10);
constant block164Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 345,10);
constant block165X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 125,10);
constant block165Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 375,10);
constant block166X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 155,10);
constant block166Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 375,10);
constant block167X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 185,10);
constant block167Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 375,10);
constant block168X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 215,10);
constant block168Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 375,10);
constant block169X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 245,10);
constant block169Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 375,10);
constant block170X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 275,10);
constant block170Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 375,10);
constant block171X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 305,10);
constant block171Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 375,10);
constant block172X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 335,10);
constant block172Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 375,10);
constant block173X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 365,10);
constant block173Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 375,10);
constant block174X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 395,10);
constant block174Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 375,10);
constant block175X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 425,10);
constant block175Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 375,10);
constant block176X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 455,10);
constant block176Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 375,10);
constant block177X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 485,10);
constant block177Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 375,10);
constant block178X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 515,10);
constant block178Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 375,10);
constant block179X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 545,10);
constant block179Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 375,10);
constant block180X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 125,10);
constant block180Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 405,10);
constant block181X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 155,10);
constant block181Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 405,10);
constant block182X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 185,10);
constant block182Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 405,10);
constant block183X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 215,10);
constant block183Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 405,10);
constant block184X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 245,10);
constant block184Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 405,10);
constant block185X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 275,10);
constant block185Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 405,10);
constant block186X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 305,10);
constant block186Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 405,10);
constant block187X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 335,10);
constant block187Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 405,10);
constant block188X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 365,10);
constant block188Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 405,10);
constant block189X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 395,10);
constant block189Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 405,10);
constant block190X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 425,10);
constant block190Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 405,10);
constant block191X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 455,10);
constant block191Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 405,10);
constant block192X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 485,10);
constant block192Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 405,10);
constant block193X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 515,10);
constant block193Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 405,10);
constant block194X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 545,10);
constant block194Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 405,10);
constant block195X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 125,10);
constant block195Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 435,10);
constant block196X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 155,10);
constant block196Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 435,10);
constant block197X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 185,10);
constant block197Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 435,10);
constant block198X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 215,10);
constant block198Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 435,10);
constant block199X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 245,10);
constant block199Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 435,10);
constant block200X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 275,10);
constant block200Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 435,10);
constant block201X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 305,10);
constant block201Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 435,10);
constant block202X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 335,10);
constant block202Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 435,10);
constant block203X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 365,10);
constant block203Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 435,10);
constant block204X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 395,10);
constant block204Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 435,10);
constant block205X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 425,10);
constant block205Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 435,10);
constant block206X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 455,10);
constant block206Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 435,10);
constant block207X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 485,10);
constant block207Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 435,10);
constant block208X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 515,10);
constant block208Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 435,10);
constant block209X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 545,10);
constant block209Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 435,10);
constant block210X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 125,10);
constant block210Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 465,10);
constant block211X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 155,10);
constant block211Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 465,10);
constant block212X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 185,10);
constant block212Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 465,10);
constant block213X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 215,10);
constant block213Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 465,10);
constant block214X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 245,10);
constant block214Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 465,10);
constant block215X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 275,10);
constant block215Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 465,10);
constant block216X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 305,10);
constant block216Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 465,10);
constant block217X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 335,10);
constant block217Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 465,10);
constant block218X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 365,10);
constant block218Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 465,10);
constant block219X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 395,10);
constant block219Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 465,10);
constant block220X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 425,10);
constant block220Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 465,10);
constant block221X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 455,10);
constant block221Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 465,10);
constant block222X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 485,10);
constant block222Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 465,10);
constant block223X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 515,10);
constant block223Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 465,10);
constant block224X : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 545,10);
constant block224Y : std_logic_vector(9 downto 0) := CONV_STD_LOGIC_VECTOR( 465,10);


begin
     chess_size <= CONV_STD_LOGIC_VECTOR(10, 10); -- assigns the chess size to be 20
get_chess_moving : process (Reset, frame_clk, state_out, button, chess_centerX, chess_centerY, chess_stepX, chess_stepY, chess_motionX, chess_motionY, counter, stop, movingX, movingY)
begin
if((state_out = "1001") or (state_out = "0001")) then
  if(Reset = '1') then   --Asynchronous Reset
      chess_motionX <= "0000000000";
      chess_motionY <= "0000000000";
      counter <= "0000000000";
      movingX <= chess_centerX;
      movingY <= chess_centerY;
  elsif(rising_edge(frame_clk)) then
    if((movingX + size >= chess_minX) and (movingX + size <= chess_maxX) and (movingY + size >= chess_minY) and (movingY + size <= chess_maxY)) then
       if(Button = x"1D") then -- move up
          if(stop = '1') then
             counter <= counter + "0000000001";
             chess_motionX <= "0000000000";
             chess_motionY <= not(chess_stepY) + '1';
          else 
             chess_motionX <= "0000000000";
             chess_motionY <= "0000000000";
          end if;
       elsif(Button = x"1B") then --  move down
          if(stop = '1') then
             counter <= counter + "0000000001";
             chess_motionX <= "0000000000";
             chess_motionY <= chess_stepY;
          else 
             chess_motionX <= "0000000000";
             chess_motionY <= "0000000000";
          end if;
       elsif(Button = x"1C") then --  move left
          if(stop = '1') then
             counter <= counter + "0000000001";
             chess_motionX <= not(chess_stepX) + '1';
             chess_motionY <= "0000000000";
          else 
             chess_motionX <= "0000000000";
             chess_motionY <= "0000000000";
          end if;
       elsif(Button = x"1C") then --  move right
          if(stop = '1') then
             counter <= counter + "0000000001";
             chess_motionX <= chess_stepX;
             chess_motionY <= "0000000000";
          else 
             chess_motionX <= "0000000000";
             chess_motionY <= "0000000000";
          end if;
       else
             chess_motionX <= chess_motionX;
             chess_motionY <= chess_motionY;
       end if;
     else
         chess_motionX <= "0000000000";
         chess_motionY <= "0000000000";
     end if;
       movingX <= movingX + chess_motionX;
       movingY <= movingY + chess_motionY;
  end if;        
 end if;
end process get_chess_moving;

get_counter_stopsig : process (counter, stop, Reset, frame_clk, state_out)
begin
    if(Reset = '1') then   --Asynchronous Reset
      counter <= "0000000000";
      stop <= '1';
    elsif(rising_edge(frame_clk)) then
      if(counter = "000001111") then -- count to 15 which the chess move 30 pixels
         stop <= '1'; 
         counter <= "000000000";
      elsif (counter = "000000000") then
         stop <= '1';
      else
         stop <= '0';
      end if;
    end if;
end process get_counter_stopsig;

stopsig <= stop;
chess_positionX <= movingX;
chess_positionY <= movingY;
chess_size <= size;

end Behavioral;


          